
module fp_multiplication_tb;

	reg [31:0] f_1;
	reg [31:0] f_2;
	wire f_nan;
	wire f_inf;
	wire [31:0] s;

	fp_multiplication uut (f_1, f_2, f_nan, f_inf, s);
	
	initial begin
			f_1 = 32'b10111101111010000100000010100001;
			f_2 = 32'b00111110110000000001000000000000;
		#5	f_1 = 32'b00111011000110100000001001110101;
			f_2 = 32'b00111101110010101100000010000011;
		#5	f_1 = 32'b00111101101001100100110000110000;
			f_2 = 32'b00111111011101000011100101011000;
		#5	$stop;
	end

endmodule
