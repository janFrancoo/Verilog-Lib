
module float_to_int_tb;

	reg [31:0] v;
	
	wire denorm;
	wire [31:0] d;
	wire p_lost;
	wire invalid;
	
	float_to_int uut (v, denorm, p_lost, invalid, d);
	
	initial begin
			v = 32'b0_10000010_10001110000101000111101; 	// 12.44
		#5	v = 32'b0_10000101_11101110001111010111000;		// 123.56
		#5	v = 32'b0_10001000_11110101000011111100111;		// 1002.123456789
		#5	v = 32'b0_11111111_00000000000000000000000;		// nan
		#5	v = 32'b0_11111111_00000100000000000000000;		// inf
		#5	v = 32'b0_11111111_00000100000000000000000;		// inf
		#5	v = 32'b1_10000001_01010000001110111001100;		// -5.25363731384
		#5	$stop;
	end

endmodule
